module GFMULT(a, b, c);
  input [3:0] a;
  input [3:0] b;
  output [3:0] c;

  assign c = ({4{b[0]}} & ((a << 0))) ^ ({4{b[1]}} & ((a << 1) ^ ({4{a[3]}} & 4'b0011))) ^ ({4{b[2]}} & ((a << 2) ^ ({4{a[3]}} & 4'b0110) ^ ({4{a[2]}} & 4'b0011))) ^ ({4{b[3]}} & ((a << 3) ^ ({4{a[3]}} & 4'b1100) ^ ({4{a[2]}} & 4'b0110) ^ ({4{a[1]}} & 4'b0011)));
endmodule
